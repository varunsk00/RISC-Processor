module register_32(out, in, clock, enable, clr);
	input [31:0] in;
	input enable;
	input clock, clr;
	output [31:0] out;

	// flip-flops
	dffe_ref flip0(out[0], in[0], clock, enable, clr);
	dffe_ref flip1(out[1], in[1], clock, enable, clr);
	dffe_ref flip2(out[2], in[2], clock, enable, clr);
	dffe_ref flip3(out[3], in[3], clock, enable, clr);
	dffe_ref flip4(out[4], in[4], clock, enable, clr);
	dffe_ref flip5(out[5], in[5], clock, enable, clr);
	dffe_ref flip6(out[6], in[6], clock, enable, clr);
	dffe_ref flip7(out[7], in[7], clock, enable, clr);
	dffe_ref flip8(out[8], in[8], clock, enable, clr);
	dffe_ref flip9(out[9], in[9], clock, enable, clr);
	dffe_ref flip10(out[10], in[10], clock, enable, clr);
	dffe_ref flip11(out[11], in[11], clock, enable, clr);
	dffe_ref flip12(out[12], in[12], clock, enable, clr);
	dffe_ref flip13(out[13], in[13], clock, enable, clr);
	dffe_ref flip14(out[14], in[14], clock, enable, clr);
	dffe_ref flip15(out[15], in[15], clock, enable, clr);
	dffe_ref flip16(out[16], in[16], clock, enable, clr);
	dffe_ref flip17(out[17], in[17], clock, enable, clr);
	dffe_ref flip18(out[18], in[18], clock, enable, clr);
	dffe_ref flip19(out[19], in[19], clock, enable, clr);
	dffe_ref flip20(out[20], in[20], clock, enable, clr);
	dffe_ref flip21(out[21], in[21], clock, enable, clr);
	dffe_ref flip22(out[22], in[22], clock, enable, clr);
	dffe_ref flip23(out[23], in[23], clock, enable, clr);
	dffe_ref flip24(out[24], in[24], clock, enable, clr);
	dffe_ref flip25(out[25], in[25], clock, enable, clr);
	dffe_ref flip26(out[26], in[26], clock, enable, clr);
	dffe_ref flip27(out[27], in[27], clock, enable, clr);
	dffe_ref flip28(out[28], in[28], clock, enable, clr);
	dffe_ref flip29(out[29], in[29], clock, enable, clr);
	dffe_ref flip30(out[30], in[30], clock, enable, clr);
	dffe_ref flip31(out[31], in[31], clock, enable, clr);
endmodule